00000093 00000113 002081B3 00000E93 00200E13 4DD19663 00100093 00100113 
002081B3 00200E93 00300E13 4BD19A63 00300093 00700113 002081B3 00A00E93 
00400E13 49D19E63 00000093 FFFF8137 002081B3 FFFF8EB7 00500E13 49D19263 
800000B7 00000113 002081B3 80000EB7 00600E13 47D19663 800000B7 FFFF8137 
002081B3 7FFF8EB7 00700E13 45D19A63 00000093 00008137 FFF10113 002081B3 
00008EB7 FFFE8E93 00800E13 43D19A63 800000B7 FFF08093 00000113 002081B3 
80000EB7 FFFE8E93 00900E13 41D19A63 800000B7 FFF08093 00008137 FFF10113 
002081B3 80008EB7 FFEE8E93 00A00E13 3FD19863 800000B7 00008137 FFF10113 
002081B3 80008EB7 FFFE8E93 00B00E13 3DD19863 800000B7 FFF08093 FFFF8137 
002081B3 7FFF8EB7 FFFE8E93 00C00E13 3BD19863 00000093 FFF00113 002081B3 
FFF00E93 00D00E13 39D19C63 FFF00093 00100113 002081B3 00000E93 00E00E13 
39D19063 FFF00093 FFF00113 002081B3 FFE00E93 00F00E13 37D19463 00100093 
80000137 FFF10113 002081B3 80000EB7 01000E13 35D19663 00D00093 00B00113 
002080B3 01800E93 01100E13 33D09A63 00E00093 00B00113 00208133 01900E93 
01200E13 31D11E63 00D00093 001080B3 01A00E93 01300E13 31D09463 00000213 
00D00093 00B00113 002081B3 00018313 00120213 00200293 FE5214E3 01800E93 
01400E13 2DD31E63 00000213 00E00093 00B00113 002081B3 00000013 00018313 
00120213 00200293 FE5212E3 01900E93 01500E13 2BD31663 00000213 00F00093 
00B00113 002081B3 00000013 00000013 00018313 00120213 00200293 FE5210E3 
01A00E93 01600E13 27D31C63 00000213 00D00093 00B00113 002081B3 00120213 
00200293 FE5216E3 01800E93 01700E13 25D19863 00000213 00E00093 00B00113 
00000013 002081B3 00120213 00200293 FE5214E3 01900E93 01800E13 23D19263 
00000213 00F00093 00B00113 00000013 00000013 002081B3 00120213 00200293 
FE5212E3 01A00E93 01900E13 1FD19A63 00000213 00D00093 00000013 00B00113 
002081B3 00120213 00200293 FE5214E3 01800E93 01A00E13 1DD19463 00000213 
00E00093 00000013 00B00113 00000013 002081B3 00120213 00200293 FE5212E3 
01900E93 01B00E13 19D19C63 00000213 00F00093 00000013 00000013 00B00113 
002081B3 00120213 00200293 FE5212E3 01A00E93 01C00E13 17D19463 00000213 
00B00113 00D00093 002081B3 00120213 00200293 FE5216E3 01800E93 01D00E13 
15D19063 00000213 00B00113 00E00093 00000013 002081B3 00120213 00200293 
FE5214E3 01900E93 01E00E13 11D19A63 00000213 00B00113 00F00093 00000013 
00000013 002081B3 00120213 00200293 FE5212E3 01A00E93 01F00E13 0FD19263 
00000213 00B00113 00000013 00D00093 002081B3 00120213 00200293 FE5214E3 
01800E93 02000E13 0BD19C63 00000213 00B00113 00000013 00E00093 00000013 
002081B3 00120213 00200293 FE5212E3 01900E93 02100E13 09D19463 00000213 
00B00113 00000013 00000013 00F00093 002081B3 00120213 00200293 FE5212E3 
01A00E93 02200E13 05D19C63 00F00093 00100133 00F00E93 02300E13 05D11263 
02000093 00008133 02000E93 02400E13 03D11863 000000B3 00000E93 02500E13 
03D09063 01000093 01E00113 00208033 00000E93 02600E13 01D01463 01C01A63 
FF000513 00000593 00B52023 FF5FF06F FF000513 00100593 00B52023 FF5FF06F 

